library ieee; 
use ieee.std_logic_1164.ALL; 
use ieee.std_logic_unsigned.ALL; 

entity pc_tb is
end pc_tb;

architecture arch of pc_tb is
begin
	process
		
	end process;
end arch;
	